
 /*
	///////////////////////////////////////////////// 
	* This part of the code taken 
	*			from LT24 Display Lab of the lecture ELEC5882
	* There is just small changing thing in this code
	* BackValue is added since when it was called firstly in top code, backValue was a need.
	* However, then design of code was changed, but it can be use in fture work.
	/////////////////////////////////////////////////
 
	* N-Bit Up Counter 
	* ---------------- 
	* By: Thomas Carpenter 
	* Date: 13/03/2017 
	* 
	* Short Description 
	* ----------------- 
	* This module is a simple up-counter with a count enable. 
	* The counter has parameter controlled width, increment, 
	* and maximum value. 
	* 
 */ 
 module UpCounterNbit #( 
	parameter WIDTH = 10, //10bit wide 
	parameter INCREMENT = 1, //Value to increment counter by each cycle 
	parameter MAX_VALUE = (2**WIDTH)-1 //Maximum value default is 2^WIDTH - 1 
 )( 
	input clock, 
	input reset, 
	input enable, //Increments when enable is high 
	input backValue, // The startin value can be different with this value(maybe it can be use for delay)
	output reg [(WIDTH-1):0] countValue //Output is declared as "WIDTH" bits wide 
 ); 
 
	always @ (posedge clock) begin 
		if (reset) begin 
			//When reset is high, set back to 0 
			countValue <= {(WIDTH){backValue}};// 1'b0}}; 
		end else if (enable) begin 
			//Otherwise counter is not in reset 
			if (countValue >= MAX_VALUE[WIDTH-1:0]) begin 
				//If the counter value is equal or exceeds the maximum value 
				countValue <= {(WIDTH){backValue}};// 1'b0}}; 
				//Reset back to 0 
			end else begin 
				//Otherwise increment 
				countValue <= countValue + INCREMENT[WIDTH-1:0]; 
			end 
		end 
	end 
 endmodule
